library IEEE;
use IEEE.std_logic_1164.all;

entity comparator_tb is
--empty
end comparator_tb;

architecture behaviour of comparator_tb is 
    component comparator is
        port(
            Ain, Bin : in STD_LOGIC;
            Gout,Sout,Eout : out STD_LOGIC
        );
    end component;

    --signal a_in, b_in, c_in, q_out, c_out: std_logic;
    signal a_in : std_logic := '0';
    signal b_in : std_logic := '0';
    signal g_out : std_ulogic;
    signal s_out : std_ulogic;
    signal e_out : std_ulogic;

    begin 
    UUT : comparator 
        port map(
            	Ain => a_in, 
            	Bin => b_in, 
            	Gout => g_out, 
            	Sout => s_out, 
            	Eout => e_out
            );

    process begin
    a_in <= '0';b_in <= '0';wait for 100 ns;
    a_in <= '0';b_in <= '1';wait for 100 ns;
    a_in <= '1';b_in <= '0';wait for 100 ns;
    a_in <= '1';b_in <= '1';wait for 100 ns;
    a_in <= '0';b_in <= '0';wait;
    end process;
end behaviour;
